// megafunction wizard: %Partial Reconfiguration v16.0%
// GENERATION: XML
// reconfig.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module reconfig (
		input  wire        clk,            //            clk.clk
		input  wire        nreset,         //         nreset.reset_n
		input  wire        pr_start,       //       pr_start.pr_start
		input  wire        double_pr,      //      double_pr.double_pr
		output wire        freeze,         //         freeze.freeze
		output wire [2:0]  status,         //         status.status
		input  wire        pr_ready_pin,   //   pr_ready_pin.pr_ready_pin
		input  wire        pr_done_pin,    //    pr_done_pin.pr_done_pin
		input  wire        pr_error_pin,   //   pr_error_pin.pr_error_pin
		input  wire        crc_error_pin,  //  crc_error_pin.crc_error_pin
		output wire        pr_request_pin, // pr_request_pin.pr_request_pin
		output wire        pr_clk_pin,     //     pr_clk_pin.pr_clk_pin
		output wire [15:0] pr_data_pin,    //    pr_data_pin.pr_data_pin
		input  wire [15:0] data,           //      avst_sink.data
		input  wire        data_valid,     //               .valid
		output wire        data_ready      //               .ready
	);

	alt_pr #(
		.PR_INTERNAL_HOST              (0),
		.ENABLE_JTAG                   (1),
		.ENABLE_AVMM_SLAVE             (0),
		.ENABLE_INTERRUPT              (0),
		.ENABLE_PRPOF_ID_CHECK         (0),
		.EXT_HOST_PRPOF_ID             (0),
		.EXT_HOST_TARGET_DEVICE_FAMILY ("Cyclone V"),
		.DATA_WIDTH_INDEX              (16),
		.CB_DATA_WIDTH                 (16),
		.ENABLE_DATA_PACKING           (1),
		.CDRATIO                       (1),
		.EDCRC_OSC_DIVIDER             (1),
		.ENABLE_ENHANCED_DECOMPRESSION (0),
		.INSTANTIATE_PR_BLOCK          (1),
		.INSTANTIATE_CRC_BLOCK         (1),
		.DEVICE_FAMILY                 ("Cyclone V")
	) reconfig_inst (
		.clk                    (clk),                  //            clk.clk
		.nreset                 (nreset),               //         nreset.reset_n
		.pr_start               (pr_start),             //       pr_start.pr_start
		.double_pr              (double_pr),            //      double_pr.double_pr
		.freeze                 (freeze),               //         freeze.freeze
		.status                 (status),               //         status.status
		.pr_ready_pin           (pr_ready_pin),         //   pr_ready_pin.pr_ready_pin
		.pr_done_pin            (pr_done_pin),          //    pr_done_pin.pr_done_pin
		.pr_error_pin           (pr_error_pin),         //   pr_error_pin.pr_error_pin
		.crc_error_pin          (crc_error_pin),        //  crc_error_pin.crc_error_pin
		.pr_request_pin         (pr_request_pin),       // pr_request_pin.pr_request_pin
		.pr_clk_pin             (pr_clk_pin),           //     pr_clk_pin.pr_clk_pin
		.pr_data_pin            (pr_data_pin),          //    pr_data_pin.pr_data_pin
		.data                   (data),                 //      avst_sink.data
		.data_valid             (data_valid),           //               .valid
		.data_ready             (data_ready),           //               .ready
		.avmm_slave_address     (1'b0),                 //    (terminated)
		.avmm_slave_read        (1'b0),                 //    (terminated)
		.avmm_slave_writedata   (16'b0000000000000000), //    (terminated)
		.avmm_slave_write       (1'b0),                 //    (terminated)
		.avmm_slave_readdata    (),                     //    (terminated)
		.avmm_slave_waitrequest (),                     //    (terminated)
		.irq                    ()                      //    (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="alt_pr" version="16.0" >
// Retrieval info: 	<generic name="PR_INTERNAL_HOST" value="false" />
// Retrieval info: 	<generic name="ENABLE_JTAG" value="true" />
// Retrieval info: 	<generic name="ENABLE_AVMM_SLAVE" value="false" />
// Retrieval info: 	<generic name="ENABLE_INTERRUPT" value="false" />
// Retrieval info: 	<generic name="ENABLE_PRPOF_ID_CHECK_UI" value="false" />
// Retrieval info: 	<generic name="EXT_HOST_PRPOF_ID" value="0" />
// Retrieval info: 	<generic name="EXT_HOST_TARGET_DEVICE_FAMILY" value="Cyclone V" />
// Retrieval info: 	<generic name="DATA_WIDTH_INDEX" value="16" />
// Retrieval info: 	<generic name="CDRATIO" value="1" />
// Retrieval info: 	<generic name="EDCRC_OSC_DIVIDER" value="1" />
// Retrieval info: 	<generic name="ENABLE_ENHANCED_DECOMPRESSION" value="false" />
// Retrieval info: 	<generic name="INSTANTIATE_PR_BLOCK" value="true" />
// Retrieval info: 	<generic name="INSTANTIATE_CRC_BLOCK" value="true" />
// Retrieval info: 	<generic name="DEVICE_FAMILY" value="Cyclone V" />
// Retrieval info: </instance>
// IPFS_FILES : reconfig.vo
// RELATED_FILES: reconfig.v, alt_pr.v, alt_pr_bitstream_host.v, alt_pr_bitstream_controller_v1.v, alt_pr_bitstream_controller_v2.v, alt_pr_cb_host.v, alt_pr_cb_interface.v, alt_pr_cb_controller_v1.v, alt_pr_cb_controller_v2.v, alt_pr_mux.sv, alt_pr_jtag_interface.v, alt_pr_width_adapter.sv, alt_pr_bitstream_compatibility_checker_int_host.v, alt_pr_bitstream_compatibility_checker_ext_host.v, alt_pr_down_converter.sv, alt_pr_fifo.sv, alt_pr_up_converter.sv, alt_pr_bitstream_decoder.sv, alt_pr_enhanced_compression_magic_words_decoder_and_suppressor.sv, alt_pr_enhanced_decompressor.sv, alt_pr_magic_fifo.sv, alt_pr_data.sv
